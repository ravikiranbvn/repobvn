module block32 ( result, cout6, cout7, cout14, cout15, cout30, cout31, a_var, b_var, var_code, anl, cin );
output [31:0] result;
input [31:0] a_var;
input [31:0] b_var;
input [3:0] var_code;
input anl, cin;
output cout6, cout7, cout14, cout15, cout30, cout31;
wire n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192;
NAND2X1 U27000 ( .A(n394), .B(n395), .Y(n496) );
NAND2X1 U27001 ( .A(n496), .B(n496), .Y(n497) );
NAND2X1 U27002 ( .A(n497), .B(n396), .Y(n233) );
NAND2X1 U271 ( .A(n233), .B(n397), .Y(n403) );
NAND2X1 U272 ( .A(b_var[15]), .B(b_var[15]), .Y(n234) );
NOR2X1 U27300 ( .A(b_var[15]), .B(n462), .Y(n498) );
NOR2X1 U27301 ( .A(n234), .B(n461), .Y(n499) );
NOR2X1 U27302 ( .A(n498), .B(n498), .Y(n500) );
NOR2X1 U27303 ( .A(n499), .B(n499), .Y(n501) );
NAND2X1 U27304 ( .A(n500), .B(n501), .Y(n235) );
NOR2X1 U27400 ( .A(b_var[15]), .B(n464), .Y(n502) );
NOR2X1 U27401 ( .A(n234), .B(n463), .Y(n503) );
NOR2X1 U27402 ( .A(n502), .B(n502), .Y(n504) );
NOR2X1 U27403 ( .A(n503), .B(n503), .Y(n505) );
NAND2X1 U27404 ( .A(n504), .B(n505), .Y(n506) );
NAND2X1 U27405 ( .A(n506), .B(n506), .Y(n507) );
NAND2X1 U27406 ( .A(n507), .B(a_var[15]), .Y(n236) );
NOR2X1 U27500 ( .A(n235), .B(a_var[15]), .Y(n508) );
NOR2X1 U27501 ( .A(n508), .B(n508), .Y(n509) );
NAND2X1 U27502 ( .A(n509), .B(n236), .Y(n326) );
NAND2X1 U27600 ( .A(anl), .B(anl), .Y(n510) );
NAND2X1 U27601 ( .A(b_var[25]), .B(b_var[25]), .Y(n511) );
NOR2X1 U27602 ( .A(n510), .B(n511), .Y(n512) );
NOR2X1 U27603 ( .A(n512), .B(n512), .Y(n513) );
NAND2X1 U27604 ( .A(n513), .B(n414), .Y(n237) );
NOR2X1 U27700 ( .A(n414), .B(n410), .Y(n514) );
NOR2X1 U27701 ( .A(n514), .B(n514), .Y(n515) );
NAND2X1 U27702 ( .A(n515), .B(n409), .Y(n516) );
NAND2X1 U27703 ( .A(n516), .B(n516), .Y(n517) );
NAND2X1 U27704 ( .A(n517), .B(n237), .Y(n417) );
NAND2X1 U278 ( .A(b_var[1]), .B(b_var[1]), .Y(n238) );
NOR2X1 U27900 ( .A(b_var[1]), .B(var_code[0]), .Y(n518) );
NOR2X1 U27901 ( .A(n238), .B(var_code[1]), .Y(n519) );
NOR2X1 U27902 ( .A(n518), .B(n518), .Y(n520) );
NOR2X1 U27903 ( .A(n519), .B(n519), .Y(n521) );
NAND2X1 U27904 ( .A(n520), .B(n521), .Y(n239) );
NOR2X1 U28000 ( .A(b_var[1]), .B(var_code[2]), .Y(n522) );
NOR2X1 U28001 ( .A(n238), .B(var_code[3]), .Y(n523) );
NOR2X1 U28002 ( .A(n522), .B(n522), .Y(n524) );
NOR2X1 U28003 ( .A(n523), .B(n523), .Y(n525) );
NAND2X1 U28004 ( .A(n524), .B(n525), .Y(n526) );
NAND2X1 U28005 ( .A(n526), .B(n526), .Y(n527) );
NAND2X1 U28006 ( .A(n527), .B(a_var[1]), .Y(n240) );
NOR2X1 U28100 ( .A(n239), .B(a_var[1]), .Y(n528) );
NOR2X1 U28101 ( .A(n528), .B(n528), .Y(n529) );
NAND2X1 U28102 ( .A(n529), .B(n240), .Y(n360) );
NAND2X1 U282 ( .A(b_var[26]), .B(b_var[26]), .Y(n241) );
NOR2X1 U28300 ( .A(b_var[26]), .B(n462), .Y(n530) );
NOR2X1 U28301 ( .A(n241), .B(n461), .Y(n531) );
NOR2X1 U28302 ( .A(n530), .B(n530), .Y(n532) );
NOR2X1 U28303 ( .A(n531), .B(n531), .Y(n533) );
NAND2X1 U28304 ( .A(n532), .B(n533), .Y(n242) );
NOR2X1 U28400 ( .A(b_var[26]), .B(n464), .Y(n534) );
NOR2X1 U28401 ( .A(n241), .B(n463), .Y(n535) );
NOR2X1 U28402 ( .A(n534), .B(n534), .Y(n536) );
NOR2X1 U28403 ( .A(n535), .B(n535), .Y(n537) );
NAND2X1 U28404 ( .A(n536), .B(n537), .Y(n538) );
NAND2X1 U28405 ( .A(n538), .B(n538), .Y(n539) );
NAND2X1 U28406 ( .A(n539), .B(a_var[26]), .Y(n243) );
NOR2X1 U28500 ( .A(n242), .B(a_var[26]), .Y(n540) );
NOR2X1 U28501 ( .A(n540), .B(n540), .Y(n541) );
NAND2X1 U28502 ( .A(n541), .B(n243), .Y(n423) );
NOR2X1 U286 ( .A(n484), .B(n483), .Y(n244) );
NOR2X1 U28700 ( .A(n287), .B(n493), .Y(n542) );
NOR2X1 U28701 ( .A(n485), .B(n244), .Y(n543) );
NOR2X1 U28702 ( .A(n542), .B(n542), .Y(n544) );
NOR2X1 U28703 ( .A(n543), .B(n543), .Y(n545) );
NOR2X1 U28704 ( .A(n544), .B(n286), .Y(n546) );
NOR2X1 U28705 ( .A(n545), .B(n482), .Y(n547) );
NOR2X1 U28706 ( .A(n546), .B(n546), .Y(n548) );
NOR2X1 U28707 ( .A(n547), .B(n547), .Y(n549) );
NAND2X1 U28708 ( .A(n548), .B(n549), .Y(cout7) );
NAND2X1 U288 ( .A(b_var[10]), .B(b_var[10]), .Y(n245) );
NOR2X1 U28900 ( .A(b_var[10]), .B(var_code[0]), .Y(n550) );
NOR2X1 U28901 ( .A(n245), .B(var_code[1]), .Y(n551) );
NOR2X1 U28902 ( .A(n550), .B(n550), .Y(n552) );
NOR2X1 U28903 ( .A(n551), .B(n551), .Y(n553) );
NAND2X1 U28904 ( .A(n552), .B(n553), .Y(n246) );
NOR2X1 U29000 ( .A(b_var[10]), .B(var_code[2]), .Y(n554) );
NOR2X1 U29001 ( .A(n245), .B(var_code[3]), .Y(n555) );
NOR2X1 U29002 ( .A(n554), .B(n554), .Y(n556) );
NOR2X1 U29003 ( .A(n555), .B(n555), .Y(n557) );
NAND2X1 U29004 ( .A(n556), .B(n557), .Y(n558) );
NAND2X1 U29005 ( .A(n558), .B(n558), .Y(n559) );
NAND2X1 U29006 ( .A(n559), .B(a_var[10]), .Y(n247) );
NOR2X1 U29100 ( .A(n246), .B(a_var[10]), .Y(n560) );
NOR2X1 U29101 ( .A(n560), .B(n560), .Y(n561) );
NAND2X1 U29102 ( .A(n561), .B(n247), .Y(n291) );
NAND2X1 U292 ( .A(b_var[11]), .B(b_var[11]), .Y(n248) );
NOR2X1 U29300 ( .A(b_var[11]), .B(var_code[0]), .Y(n562) );
NOR2X1 U29301 ( .A(n248), .B(var_code[1]), .Y(n563) );
NOR2X1 U29302 ( .A(n562), .B(n562), .Y(n564) );
NOR2X1 U29303 ( .A(n563), .B(n563), .Y(n565) );
NAND2X1 U29304 ( .A(n564), .B(n565), .Y(n249) );
NOR2X1 U29400 ( .A(b_var[11]), .B(var_code[2]), .Y(n566) );
NOR2X1 U29401 ( .A(n248), .B(var_code[3]), .Y(n567) );
NOR2X1 U29402 ( .A(n566), .B(n566), .Y(n568) );
NOR2X1 U29403 ( .A(n567), .B(n567), .Y(n569) );
NAND2X1 U29404 ( .A(n568), .B(n569), .Y(n570) );
NAND2X1 U29405 ( .A(n570), .B(n570), .Y(n571) );
NAND2X1 U29406 ( .A(n571), .B(a_var[11]), .Y(n250) );
NOR2X1 U29500 ( .A(n249), .B(a_var[11]), .Y(n572) );
NOR2X1 U29501 ( .A(n572), .B(n572), .Y(n573) );
NAND2X1 U29502 ( .A(n573), .B(n250), .Y(n296) );
NOR2X1 U29600 ( .A(cin), .B(n495), .Y(n574) );
NOR2X1 U29601 ( .A(n574), .B(n574), .Y(n575) );
NAND2X1 U29602 ( .A(n575), .B(n359), .Y(n251) );
NOR2X1 U29700 ( .A(n360), .B(n251), .Y(n576) );
NOR2X1 U29701 ( .A(n360), .B(n576), .Y(n577) );
NOR2X1 U29702 ( .A(n576), .B(n251), .Y(n578) );
NOR2X1 U29703 ( .A(n577), .B(n578), .Y(result[1]) );
NAND2X1 U29800 ( .A(n349), .B(n339), .Y(n579) );
NAND2X1 U29801 ( .A(n336), .B(n339), .Y(n580) );
NAND2X1 U29802 ( .A(n579), .B(n579), .Y(n581) );
NAND2X1 U29803 ( .A(n580), .B(n580), .Y(n582) );
NAND2X1 U29804 ( .A(n581), .B(n350), .Y(n583) );
NAND2X1 U29805 ( .A(n583), .B(n583), .Y(n584) );
NOR2X1 U29806 ( .A(n584), .B(n582), .Y(result[17]) );
NOR2X1 U29900 ( .A(n400), .B(n403), .Y(n585) );
NOR2X1 U29901 ( .A(n585), .B(n585), .Y(n586) );
NAND2X1 U29902 ( .A(n586), .B(n405), .Y(n252) );
NOR2X1 U30000 ( .A(n406), .B(n252), .Y(n587) );
NOR2X1 U30001 ( .A(n406), .B(n587), .Y(n588) );
NOR2X1 U30002 ( .A(n587), .B(n252), .Y(n589) );
NOR2X1 U30003 ( .A(n588), .B(n589), .Y(result[24]) );
NAND2X1 U30100 ( .A(n448), .B(n435), .Y(n590) );
NAND2X1 U30101 ( .A(n432), .B(n435), .Y(n591) );
NAND2X1 U30102 ( .A(n590), .B(n590), .Y(n592) );
NAND2X1 U30103 ( .A(n591), .B(n591), .Y(n593) );
NAND2X1 U30104 ( .A(n592), .B(n449), .Y(n594) );
NAND2X1 U30105 ( .A(n594), .B(n594), .Y(n595) );
NOR2X1 U30106 ( .A(n595), .B(n593), .Y(result[28]) );
NOR2X1 U30200 ( .A(n494), .B(n493), .Y(n596) );
NOR2X1 U30201 ( .A(n491), .B(n490), .Y(n597) );
NOR2X1 U30202 ( .A(n596), .B(n596), .Y(n598) );
NOR2X1 U30203 ( .A(n597), .B(n597), .Y(n599) );
NOR2X1 U30204 ( .A(n598), .B(n492), .Y(n600) );
NOR2X1 U30205 ( .A(n600), .B(n600), .Y(n601) );
NAND2X1 U30206 ( .A(n601), .B(n599), .Y(cout31) );
NAND2X1 U303 ( .A(n457), .B(n457), .Y(result[30]) );
NOR2X1 U30400 ( .A(n440), .B(n455), .Y(n602) );
NOR2X1 U30401 ( .A(n602), .B(n602), .Y(n603) );
NAND2X1 U30402 ( .A(n603), .B(n439), .Y(result[29]) );
NAND2X1 U305 ( .A(n440), .B(n455), .Y(n439) );
NAND2X1 U306 ( .A(n435), .B(n434), .Y(n440) );
NOR2X1 U30700 ( .A(n431), .B(n429), .Y(n604) );
NOR2X1 U30701 ( .A(n604), .B(n604), .Y(n605) );
NOR2X1 U30702 ( .A(n605), .B(n428), .Y(n606) );
NOR2X1 U30703 ( .A(n606), .B(n606), .Y(n607) );
NAND2X1 U30704 ( .A(n607), .B(n424), .Y(result[27]) );
NAND2X1 U308 ( .A(n416), .B(n423), .Y(n415) );
NAND2X1 U309 ( .A(n417), .B(n422), .Y(n416) );
NAND2X1 U310 ( .A(n414), .B(n414), .Y(n408) );
NOR2X1 U31100 ( .A(n389), .B(n396), .Y(n608) );
NOR2X1 U31101 ( .A(n608), .B(n608), .Y(n609) );
NAND2X1 U31102 ( .A(n609), .B(n388), .Y(result[23]) );
NAND2X1 U312 ( .A(n389), .B(n396), .Y(n388) );
NOR2X1 U31300 ( .A(n379), .B(n409), .Y(n610) );
NOR2X1 U31301 ( .A(n610), .B(n610), .Y(n611) );
NAND2X1 U31302 ( .A(n611), .B(n381), .Y(n380) );
NAND2X1 U314 ( .A(n409), .B(n409), .Y(n400) );
NAND2X1 U315 ( .A(n368), .B(n368), .Y(result[20]) );
NAND2X1 U316 ( .A(n358), .B(n358), .Y(result[19]) );
NOR2X1 U31700 ( .A(n344), .B(n356), .Y(n612) );
NOR2X1 U31701 ( .A(n612), .B(n612), .Y(n613) );
NAND2X1 U31702 ( .A(n613), .B(n343), .Y(result[18]) );
NAND2X1 U318 ( .A(n344), .B(n356), .Y(n343) );
NAND2X1 U319 ( .A(n339), .B(n338), .Y(n344) );
NOR2X1 U32000 ( .A(n333), .B(n333), .Y(n614) );
NOR2X1 U32001 ( .A(cout15), .B(cout15), .Y(n615) );
NOR2X1 U32002 ( .A(n614), .B(n615), .Y(n616) );
NOR2X1 U32003 ( .A(n333), .B(cout15), .Y(n617) );
NOR2X1 U32004 ( .A(n616), .B(n616), .Y(n618) );
NOR2X1 U32005 ( .A(n617), .B(n617), .Y(n619) );
NAND2X1 U32006 ( .A(n618), .B(n619), .Y(result[16]) );
NOR2X1 U32100 ( .A(n326), .B(n326), .Y(n620) );
NOR2X1 U32101 ( .A(cout14), .B(cout14), .Y(n621) );
NOR2X1 U32102 ( .A(n620), .B(n621), .Y(n622) );
NOR2X1 U32103 ( .A(n326), .B(cout14), .Y(n623) );
NOR2X1 U32104 ( .A(n622), .B(n622), .Y(n624) );
NOR2X1 U32105 ( .A(n623), .B(n623), .Y(n625) );
NAND2X1 U32106 ( .A(n624), .B(n625), .Y(result[15]) );
NAND2X1 U322 ( .A(n316), .B(n322), .Y(n315) );
NOR2X1 U32300 ( .A(a_var[31]), .B(n466), .Y(n626) );
NOR2X1 U32301 ( .A(n626), .B(n626), .Y(n627) );
NAND2X1 U32302 ( .A(n627), .B(n465), .Y(n490) );
NAND2X1 U324 ( .A(cout30), .B(cout30), .Y(n491) );
NOR2X1 U32500 ( .A(n306), .B(n306), .Y(n628) );
NOR2X1 U32501 ( .A(n307), .B(n307), .Y(n629) );
NOR2X1 U32502 ( .A(n628), .B(n629), .Y(n630) );
NOR2X1 U32503 ( .A(n306), .B(n307), .Y(n631) );
NOR2X1 U32504 ( .A(n630), .B(n630), .Y(n632) );
NOR2X1 U32505 ( .A(n631), .B(n631), .Y(n633) );
NAND2X1 U32506 ( .A(n632), .B(n633), .Y(result[12]) );
NOR2X1 U32600 ( .A(n291), .B(n290), .Y(n634) );
NOR2X1 U32601 ( .A(n634), .B(n634), .Y(n635) );
NAND2X1 U32602 ( .A(n635), .B(n292), .Y(result[10]) );
NAND2X1 U32700 ( .A(n489), .B(n488), .Y(n636) );
NAND2X1 U32701 ( .A(n636), .B(n636), .Y(n637) );
NOR2X1 U32702 ( .A(n637), .B(n487), .Y(result[9]) );
NOR2X1 U32800 ( .A(cout7), .B(cout7), .Y(n638) );
NOR2X1 U32801 ( .A(n486), .B(n486), .Y(n639) );
NOR2X1 U32802 ( .A(n638), .B(n639), .Y(n640) );
NOR2X1 U32803 ( .A(cout7), .B(n486), .Y(n641) );
NOR2X1 U32804 ( .A(n640), .B(n640), .Y(n642) );
NOR2X1 U32805 ( .A(n641), .B(n641), .Y(n643) );
NAND2X1 U32806 ( .A(n642), .B(n643), .Y(result[8]) );
NAND2X1 U329 ( .A(n477), .B(n476), .Y(n479) );
NAND2X1 U33000 ( .A(n477), .B(n475), .Y(n644) );
NAND2X1 U33001 ( .A(n644), .B(n644), .Y(n645) );
NAND2X1 U33002 ( .A(n645), .B(n478), .Y(n646) );
NAND2X1 U33003 ( .A(n646), .B(n646), .Y(n647) );
NOR2X1 U33004 ( .A(n647), .B(n474), .Y(n480) );
NAND2X1 U331 ( .A(n475), .B(n475), .Y(n476) );
NAND2X1 U33200 ( .A(n472), .B(n471), .Y(n648) );
NAND2X1 U33201 ( .A(n648), .B(n648), .Y(n649) );
NOR2X1 U33202 ( .A(n649), .B(n470), .Y(result[4]) );
NAND2X1 U33300 ( .A(n469), .B(n468), .Y(n650) );
NAND2X1 U33301 ( .A(n650), .B(n650), .Y(n651) );
NOR2X1 U33302 ( .A(n651), .B(n467), .Y(result[3]) );
NOR2X1 U33400 ( .A(n443), .B(n442), .Y(n652) );
NOR2X1 U33401 ( .A(n652), .B(n652), .Y(n653) );
NAND2X1 U33402 ( .A(n653), .B(n441), .Y(result[2]) );
NOR2X1 U33500 ( .A(n495), .B(n495), .Y(n654) );
NOR2X1 U33501 ( .A(cin), .B(cin), .Y(n655) );
NOR2X1 U33502 ( .A(n654), .B(n655), .Y(n656) );
NOR2X1 U33503 ( .A(n495), .B(cin), .Y(n657) );
NOR2X1 U33504 ( .A(n656), .B(n656), .Y(n658) );
NOR2X1 U33505 ( .A(n657), .B(n657), .Y(n659) );
NAND2X1 U33506 ( .A(n658), .B(n659), .Y(result[0]) );
NOR2X1 U33600 ( .A(n455), .B(n454), .Y(n660) );
NOR2X1 U33601 ( .A(n660), .B(n660), .Y(n661) );
NAND2X1 U33602 ( .A(n661), .B(n453), .Y(n456) );
NAND2X1 U337 ( .A(n431), .B(n430), .Y(n449) );
NAND2X1 U338 ( .A(n374), .B(n367), .Y(n372) );
NAND2X1 U339 ( .A(n366), .B(n357), .Y(n364) );
NAND2X1 U340 ( .A(n335), .B(n334), .Y(n350) );
NOR2X1 U34100 ( .A(n309), .B(n308), .Y(n662) );
NOR2X1 U34101 ( .A(n662), .B(n662), .Y(n663) );
NOR2X1 U34102 ( .A(n663), .B(n307), .Y(n321) );
NAND2X1 U342 ( .A(n477), .B(n477), .Y(n473) );
NOR2X1 U34300 ( .A(a_var[2]), .B(n283), .Y(n664) );
NOR2X1 U34301 ( .A(n664), .B(n664), .Y(n665) );
NAND2X1 U34302 ( .A(n665), .B(n282), .Y(n442) );
NAND2X1 U34400 ( .A(b_var[0]), .B(b_var[0]), .Y(n666) );
NAND2X1 U34401 ( .A(n495), .B(n495), .Y(n667) );
NOR2X1 U34402 ( .A(n666), .B(n667), .Y(n668) );
NOR2X1 U34403 ( .A(n668), .B(n668), .Y(n669) );
NAND2X1 U34404 ( .A(n669), .B(n360), .Y(n278) );
NOR2X1 U34500 ( .A(n277), .B(n493), .Y(n670) );
NOR2X1 U34501 ( .A(n670), .B(n670), .Y(n671) );
NAND2X1 U34502 ( .A(n671), .B(n495), .Y(n359) );
NOR2X1 U34600 ( .A(a_var[0]), .B(n276), .Y(n672) );
NOR2X1 U34601 ( .A(n672), .B(n672), .Y(n673) );
NAND2X1 U34602 ( .A(n673), .B(n275), .Y(n495) );
NOR2X1 U34700 ( .A(a_var[3]), .B(n274), .Y(n674) );
NOR2X1 U34701 ( .A(n674), .B(n674), .Y(n675) );
NAND2X1 U34702 ( .A(n675), .B(n273), .Y(n468) );
NOR2X1 U34800 ( .A(a_var[4]), .B(n271), .Y(n676) );
NOR2X1 U34801 ( .A(n676), .B(n676), .Y(n677) );
NAND2X1 U34802 ( .A(n677), .B(n270), .Y(n471) );
NOR2X1 U34900 ( .A(a_var[5]), .B(n266), .Y(n678) );
NOR2X1 U34901 ( .A(n265), .B(n264), .Y(n679) );
NOR2X1 U34902 ( .A(n678), .B(n678), .Y(n680) );
NOR2X1 U34903 ( .A(n679), .B(n679), .Y(n681) );
NAND2X1 U34904 ( .A(n680), .B(n681), .Y(n477) );
NOR2X1 U35000 ( .A(a_var[6]), .B(n263), .Y(n682) );
NOR2X1 U35001 ( .A(n262), .B(n261), .Y(n683) );
NOR2X1 U35002 ( .A(n682), .B(n682), .Y(n684) );
NOR2X1 U35003 ( .A(n683), .B(n683), .Y(n685) );
NAND2X1 U35004 ( .A(n684), .B(n685), .Y(n284) );
NOR2X1 U35100 ( .A(a_var[7]), .B(n260), .Y(n686) );
NOR2X1 U35101 ( .A(n259), .B(n258), .Y(n687) );
NOR2X1 U35102 ( .A(n686), .B(n686), .Y(n688) );
NOR2X1 U35103 ( .A(n687), .B(n687), .Y(n689) );
NAND2X1 U35104 ( .A(n688), .B(n689), .Y(n287) );
NOR2X1 U35200 ( .A(b_var[7]), .B(var_code[2]), .Y(n690) );
NOR2X1 U35201 ( .A(n286), .B(var_code[3]), .Y(n691) );
NOR2X1 U35202 ( .A(n690), .B(n690), .Y(n692) );
NOR2X1 U35203 ( .A(n691), .B(n691), .Y(n693) );
NAND2X1 U35204 ( .A(n692), .B(n693), .Y(n258) );
NOR2X1 U35300 ( .A(b_var[7]), .B(var_code[0]), .Y(n694) );
NOR2X1 U35301 ( .A(n286), .B(var_code[1]), .Y(n695) );
NOR2X1 U35302 ( .A(n694), .B(n694), .Y(n696) );
NOR2X1 U35303 ( .A(n695), .B(n695), .Y(n697) );
NAND2X1 U35304 ( .A(n696), .B(n697), .Y(n260) );
NOR2X1 U35400 ( .A(a_var[8]), .B(n257), .Y(n698) );
NOR2X1 U35401 ( .A(n698), .B(n698), .Y(n699) );
NAND2X1 U35402 ( .A(n699), .B(n256), .Y(n486) );
NOR2X1 U35500 ( .A(b_var[8]), .B(n462), .Y(n700) );
NOR2X1 U35501 ( .A(n288), .B(n461), .Y(n701) );
NOR2X1 U35502 ( .A(n700), .B(n700), .Y(n702) );
NOR2X1 U35503 ( .A(n701), .B(n701), .Y(n703) );
NAND2X1 U35504 ( .A(n702), .B(n703), .Y(n257) );
NOR2X1 U35600 ( .A(a_var[9]), .B(n255), .Y(n704) );
NOR2X1 U35601 ( .A(n704), .B(n704), .Y(n705) );
NAND2X1 U35602 ( .A(n705), .B(n254), .Y(n488) );
NAND2X1 U357 ( .A(n312), .B(n312), .Y(n302) );
NOR2X1 U35800 ( .A(n326), .B(n325), .Y(n706) );
NOR2X1 U35801 ( .A(n706), .B(n706), .Y(n707) );
NAND2X1 U35802 ( .A(n707), .B(n324), .Y(n332) );
NOR2X1 U35900 ( .A(n320), .B(n319), .Y(n708) );
NOR2X1 U35901 ( .A(n708), .B(n708), .Y(n709) );
NAND2X1 U35902 ( .A(n709), .B(n318), .Y(n325) );
NOR2X1 U36000 ( .A(a_var[14]), .B(n314), .Y(n710) );
NOR2X1 U36001 ( .A(n710), .B(n710), .Y(n711) );
NAND2X1 U36002 ( .A(n711), .B(n313), .Y(n319) );
NOR2X1 U36100 ( .A(b_var[14]), .B(n462), .Y(n712) );
NOR2X1 U36101 ( .A(n317), .B(n461), .Y(n713) );
NOR2X1 U36102 ( .A(n712), .B(n712), .Y(n714) );
NOR2X1 U36103 ( .A(n713), .B(n713), .Y(n715) );
NAND2X1 U36104 ( .A(n714), .B(n715), .Y(n314) );
NOR2X1 U36200 ( .A(a_var[12]), .B(n295), .Y(n716) );
NOR2X1 U36201 ( .A(n716), .B(n716), .Y(n717) );
NAND2X1 U36202 ( .A(n717), .B(n294), .Y(n300) );
NOR2X1 U36300 ( .A(b_var[12]), .B(n462), .Y(n718) );
NOR2X1 U36301 ( .A(n304), .B(n461), .Y(n719) );
NOR2X1 U36302 ( .A(n718), .B(n718), .Y(n720) );
NOR2X1 U36303 ( .A(n719), .B(n719), .Y(n721) );
NAND2X1 U36304 ( .A(n720), .B(n721), .Y(n295) );
NOR2X1 U36400 ( .A(a_var[13]), .B(n299), .Y(n722) );
NOR2X1 U36401 ( .A(n722), .B(n722), .Y(n723) );
NAND2X1 U36402 ( .A(n723), .B(n298), .Y(n312) );
NOR2X1 U36500 ( .A(b_var[13]), .B(n462), .Y(n724) );
NOR2X1 U36501 ( .A(n303), .B(n461), .Y(n725) );
NOR2X1 U36502 ( .A(n724), .B(n724), .Y(n726) );
NOR2X1 U36503 ( .A(n725), .B(n725), .Y(n727) );
NAND2X1 U36504 ( .A(n726), .B(n727), .Y(n299) );
NOR2X1 U36600 ( .A(a_var[16]), .B(n328), .Y(n728) );
NOR2X1 U36601 ( .A(n728), .B(n728), .Y(n729) );
NAND2X1 U36602 ( .A(n729), .B(n327), .Y(n333) );
NOR2X1 U36700 ( .A(a_var[17]), .B(n330), .Y(n730) );
NOR2X1 U36701 ( .A(n730), .B(n730), .Y(n731) );
NAND2X1 U36702 ( .A(n731), .B(n329), .Y(n351) );
NOR2X1 U36800 ( .A(a_var[18]), .B(n342), .Y(n732) );
NOR2X1 U36801 ( .A(n732), .B(n732), .Y(n733) );
NAND2X1 U36802 ( .A(n733), .B(n341), .Y(n356) );
NOR2X1 U36900 ( .A(a_var[19]), .B(n347), .Y(n734) );
NOR2X1 U36901 ( .A(n346), .B(n345), .Y(n735) );
NOR2X1 U36902 ( .A(n734), .B(n734), .Y(n736) );
NOR2X1 U36903 ( .A(n735), .B(n735), .Y(n737) );
NAND2X1 U36904 ( .A(n736), .B(n737), .Y(n366) );
NOR2X1 U37000 ( .A(a_var[20]), .B(n363), .Y(n738) );
NOR2X1 U37001 ( .A(n362), .B(n361), .Y(n739) );
NOR2X1 U37002 ( .A(n738), .B(n738), .Y(n740) );
NOR2X1 U37003 ( .A(n739), .B(n739), .Y(n741) );
NAND2X1 U37004 ( .A(n740), .B(n741), .Y(n374) );
NOR2X1 U37100 ( .A(n423), .B(n422), .Y(n742) );
NOR2X1 U37101 ( .A(n742), .B(n742), .Y(n743) );
NAND2X1 U37102 ( .A(n743), .B(n421), .Y(n428) );
NAND2X1 U372 ( .A(n382), .B(n382), .Y(n383) );
NAND2X1 U373 ( .A(n382), .B(n381), .Y(n394) );
NOR2X1 U37400 ( .A(n378), .B(n493), .Y(n744) );
NOR2X1 U37401 ( .A(n744), .B(n744), .Y(n745) );
NAND2X1 U37402 ( .A(n745), .B(n379), .Y(n381) );
NOR2X1 U37500 ( .A(a_var[22]), .B(n377), .Y(n746) );
NOR2X1 U37501 ( .A(n746), .B(n746), .Y(n747) );
NAND2X1 U37502 ( .A(n747), .B(n376), .Y(n382) );
NOR2X1 U37600 ( .A(b_var[22]), .B(var_code[0]), .Y(n748) );
NOR2X1 U37601 ( .A(n375), .B(var_code[1]), .Y(n749) );
NOR2X1 U37602 ( .A(n748), .B(n748), .Y(n750) );
NOR2X1 U37603 ( .A(n749), .B(n749), .Y(n751) );
NAND2X1 U37604 ( .A(n750), .B(n751), .Y(n377) );
NOR2X1 U37700 ( .A(a_var[21]), .B(n371), .Y(n752) );
NOR2X1 U37701 ( .A(n370), .B(n369), .Y(n753) );
NOR2X1 U37702 ( .A(n752), .B(n752), .Y(n754) );
NOR2X1 U37703 ( .A(n753), .B(n753), .Y(n755) );
NAND2X1 U37704 ( .A(n754), .B(n755), .Y(n384) );
NOR2X1 U37800 ( .A(a_var[23]), .B(n387), .Y(n756) );
NOR2X1 U37801 ( .A(n386), .B(n385), .Y(n757) );
NOR2X1 U37802 ( .A(n756), .B(n756), .Y(n758) );
NOR2X1 U37803 ( .A(n757), .B(n757), .Y(n759) );
NAND2X1 U37804 ( .A(n758), .B(n759), .Y(n399) );
NOR2X1 U37900 ( .A(a_var[24]), .B(n392), .Y(n760) );
NOR2X1 U37901 ( .A(n760), .B(n760), .Y(n761) );
NAND2X1 U37902 ( .A(n761), .B(n391), .Y(n406) );
NOR2X1 U38000 ( .A(b_var[24]), .B(n462), .Y(n762) );
NOR2X1 U38001 ( .A(n390), .B(n461), .Y(n763) );
NOR2X1 U38002 ( .A(n762), .B(n762), .Y(n764) );
NOR2X1 U38003 ( .A(n763), .B(n763), .Y(n765) );
NAND2X1 U38004 ( .A(n764), .B(n765), .Y(n392) );
NOR2X1 U38100 ( .A(a_var[25]), .B(n402), .Y(n766) );
NOR2X1 U38101 ( .A(n766), .B(n766), .Y(n767) );
NAND2X1 U38102 ( .A(n767), .B(n401), .Y(n414) );
NOR2X1 U38200 ( .A(b_var[25]), .B(n462), .Y(n768) );
NOR2X1 U38201 ( .A(n411), .B(n461), .Y(n769) );
NOR2X1 U38202 ( .A(n768), .B(n768), .Y(n770) );
NOR2X1 U38203 ( .A(n769), .B(n769), .Y(n771) );
NAND2X1 U38204 ( .A(n770), .B(n771), .Y(n402) );
NOR2X1 U38300 ( .A(a_var[27]), .B(n420), .Y(n772) );
NOR2X1 U38301 ( .A(n419), .B(n418), .Y(n773) );
NOR2X1 U38302 ( .A(n772), .B(n772), .Y(n774) );
NOR2X1 U38303 ( .A(n773), .B(n773), .Y(n775) );
NAND2X1 U38304 ( .A(n774), .B(n775), .Y(n429) );
NOR2X1 U38400 ( .A(a_var[28]), .B(n426), .Y(n776) );
NOR2X1 U38401 ( .A(n776), .B(n776), .Y(n777) );
NAND2X1 U38402 ( .A(n777), .B(n425), .Y(n450) );
NAND2X1 U385 ( .A(var_code[3]), .B(var_code[3]), .Y(n463) );
NAND2X1 U386 ( .A(var_code[2]), .B(var_code[2]), .Y(n464) );
NAND2X1 U387 ( .A(var_code[1]), .B(var_code[1]), .Y(n461) );
NAND2X1 U388 ( .A(var_code[0]), .B(var_code[0]), .Y(n462) );
NOR2X1 U38900 ( .A(a_var[29]), .B(n438), .Y(n778) );
NOR2X1 U38901 ( .A(n778), .B(n778), .Y(n779) );
NAND2X1 U38902 ( .A(n779), .B(n437), .Y(n455) );
NAND2X1 U390 ( .A(anl), .B(anl), .Y(n493) );
NOR2X1 U39100 ( .A(a_var[30]), .B(n446), .Y(n780) );
NOR2X1 U39101 ( .A(n445), .B(n444), .Y(n781) );
NOR2X1 U39102 ( .A(n780), .B(n780), .Y(n782) );
NOR2X1 U39103 ( .A(n781), .B(n781), .Y(n783) );
NAND2X1 U39104 ( .A(n782), .B(n783), .Y(n460) );
NAND2X1 U392 ( .A(n450), .B(n450), .Y(n432) );
NAND2X1 U39300 ( .A(n410), .B(n409), .Y(n784) );
NAND2X1 U39301 ( .A(n784), .B(n784), .Y(n785) );
NOR2X1 U39302 ( .A(n785), .B(n413), .Y(n407) );
NAND2X1 U39400 ( .A(n394), .B(n394), .Y(n786) );
NAND2X1 U39401 ( .A(n400), .B(n400), .Y(n787) );
NAND2X1 U39402 ( .A(n786), .B(n787), .Y(n788) );
NOR2X1 U39403 ( .A(n789), .B(n398), .Y(n389) );
NAND2X1 U39404 ( .A(n788), .B(n788), .Y(n789) );
NAND2X1 U395 ( .A(n351), .B(n351), .Y(n336) );
NAND2X1 U396 ( .A(n490), .B(n490), .Y(n494) );
NOR2X1 U39700 ( .A(b_var[31]), .B(n464), .Y(n790) );
NOR2X1 U39701 ( .A(n492), .B(n463), .Y(n791) );
NOR2X1 U39702 ( .A(n790), .B(n790), .Y(n792) );
NOR2X1 U39703 ( .A(n791), .B(n791), .Y(n793) );
NAND2X1 U39704 ( .A(n792), .B(n793), .Y(n794) );
NAND2X1 U39705 ( .A(n794), .B(n794), .Y(n795) );
NAND2X1 U39706 ( .A(n795), .B(a_var[31]), .Y(n465) );
NAND2X1 U398 ( .A(b_var[31]), .B(b_var[31]), .Y(n492) );
NOR2X1 U39900 ( .A(n485), .B(n485), .Y(n796) );
NOR2X1 U39901 ( .A(cout6), .B(cout6), .Y(n797) );
NOR2X1 U39902 ( .A(n796), .B(n797), .Y(n798) );
NOR2X1 U39903 ( .A(n485), .B(cout6), .Y(n799) );
NOR2X1 U39904 ( .A(n798), .B(n798), .Y(n800) );
NOR2X1 U39905 ( .A(n799), .B(n799), .Y(n801) );
NAND2X1 U39906 ( .A(n800), .B(n801), .Y(result[7]) );
NAND2X1 U40000 ( .A(n481), .B(n480), .Y(n802) );
NAND2X1 U40001 ( .A(n478), .B(n480), .Y(n803) );
NAND2X1 U40002 ( .A(n802), .B(n802), .Y(n804) );
NAND2X1 U40003 ( .A(n803), .B(n803), .Y(n805) );
NAND2X1 U40004 ( .A(n804), .B(n479), .Y(n806) );
NAND2X1 U40005 ( .A(n806), .B(n806), .Y(n807) );
NOR2X1 U40006 ( .A(n807), .B(n805), .Y(result[6]) );
NAND2X1 U40100 ( .A(n484), .B(n484), .Y(n808) );
NAND2X1 U40101 ( .A(n483), .B(n483), .Y(n809) );
NAND2X1 U40102 ( .A(n808), .B(n809), .Y(n810) );
NOR2X1 U40103 ( .A(n811), .B(n482), .Y(cout6) );
NAND2X1 U40104 ( .A(n810), .B(n810), .Y(n811) );
NAND2X1 U402 ( .A(n325), .B(n323), .Y(cout14) );
NOR2X1 U40300 ( .A(n335), .B(n332), .Y(n812) );
NOR2X1 U40301 ( .A(n812), .B(n812), .Y(cout15) );
NOR2X1 U40400 ( .A(n460), .B(n459), .Y(n813) );
NOR2X1 U40401 ( .A(n813), .B(n813), .Y(n814) );
NOR2X1 U40402 ( .A(n814), .B(n493), .Y(n815) );
NOR2X1 U40403 ( .A(n815), .B(n815), .Y(n816) );
NAND2X1 U40404 ( .A(n816), .B(n458), .Y(cout30) );
NAND2X1 U405 ( .A(n460), .B(n456), .Y(n458) );
NOR2X1 U40600 ( .A(n374), .B(n373), .Y(n817) );
NOR2X1 U40601 ( .A(n817), .B(n817), .Y(n818) );
NOR2X1 U40602 ( .A(n818), .B(n493), .Y(n819) );
NOR2X1 U40603 ( .A(n819), .B(n819), .Y(n820) );
NAND2X1 U40604 ( .A(n820), .B(n372), .Y(n409) );
NOR2X1 U40700 ( .A(n366), .B(n365), .Y(n821) );
NOR2X1 U40701 ( .A(n821), .B(n821), .Y(n822) );
NOR2X1 U40702 ( .A(n822), .B(n493), .Y(n823) );
NOR2X1 U40703 ( .A(n823), .B(n823), .Y(n824) );
NAND2X1 U40704 ( .A(n824), .B(n364), .Y(n367) );
NAND2X1 U408 ( .A(n322), .B(n321), .Y(n323) );
NAND2X1 U40900 ( .A(b_var[11]), .B(n297), .Y(n825) );
NAND2X1 U40901 ( .A(n296), .B(n297), .Y(n826) );
NAND2X1 U40902 ( .A(n825), .B(n825), .Y(n827) );
NAND2X1 U40903 ( .A(n826), .B(n826), .Y(n828) );
NAND2X1 U40904 ( .A(n827), .B(anl), .Y(n829) );
NAND2X1 U40905 ( .A(n829), .B(n829), .Y(n830) );
NOR2X1 U40906 ( .A(n830), .B(n828), .Y(n307) );
NAND2X1 U410 ( .A(n296), .B(n293), .Y(n297) );
NAND2X1 U41100 ( .A(b_var[10]), .B(n292), .Y(n831) );
NAND2X1 U41101 ( .A(n291), .B(n292), .Y(n832) );
NAND2X1 U41102 ( .A(n831), .B(n831), .Y(n833) );
NAND2X1 U41103 ( .A(n832), .B(n832), .Y(n834) );
NAND2X1 U41104 ( .A(n833), .B(anl), .Y(n835) );
NAND2X1 U41105 ( .A(n835), .B(n835), .Y(n836) );
NOR2X1 U41106 ( .A(n836), .B(n834), .Y(n293) );
NAND2X1 U412 ( .A(n291), .B(n290), .Y(n292) );
NAND2X1 U41300 ( .A(b_var[9]), .B(anl), .Y(n837) );
NAND2X1 U41301 ( .A(n837), .B(n837), .Y(n838) );
NAND2X1 U41302 ( .A(n838), .B(n488), .Y(n839) );
NAND2X1 U41303 ( .A(n839), .B(n839), .Y(n840) );
NOR2X1 U41304 ( .A(n840), .B(n487), .Y(n290) );
NAND2X1 U414 ( .A(n287), .B(n287), .Y(n485) );
NAND2X1 U41500 ( .A(n493), .B(n493), .Y(n841) );
NAND2X1 U41501 ( .A(n285), .B(n285), .Y(n842) );
NAND2X1 U41502 ( .A(n841), .B(n842), .Y(n843) );
NOR2X1 U41503 ( .A(n844), .B(n478), .Y(n482) );
NAND2X1 U41504 ( .A(n843), .B(n843), .Y(n844) );
NAND2X1 U416 ( .A(n478), .B(n481), .Y(n483) );
NAND2X1 U417 ( .A(n284), .B(n284), .Y(n478) );
NAND2X1 U41800 ( .A(b_var[4]), .B(anl), .Y(n845) );
NAND2X1 U41801 ( .A(n845), .B(n845), .Y(n846) );
NAND2X1 U41802 ( .A(n846), .B(n471), .Y(n847) );
NAND2X1 U41803 ( .A(n847), .B(n847), .Y(n848) );
NOR2X1 U41804 ( .A(n848), .B(n470), .Y(n475) );
NAND2X1 U41900 ( .A(b_var[3]), .B(anl), .Y(n849) );
NAND2X1 U41901 ( .A(n849), .B(n849), .Y(n850) );
NAND2X1 U41902 ( .A(n850), .B(n468), .Y(n851) );
NAND2X1 U41903 ( .A(n851), .B(n851), .Y(n852) );
NOR2X1 U41904 ( .A(n852), .B(n467), .Y(n472) );
NAND2X1 U42000 ( .A(b_var[2]), .B(n441), .Y(n853) );
NAND2X1 U42001 ( .A(n442), .B(n441), .Y(n854) );
NAND2X1 U42002 ( .A(n853), .B(n853), .Y(n855) );
NAND2X1 U42003 ( .A(n854), .B(n854), .Y(n856) );
NAND2X1 U42004 ( .A(n855), .B(anl), .Y(n857) );
NAND2X1 U42005 ( .A(n857), .B(n857), .Y(n858) );
NOR2X1 U42006 ( .A(n858), .B(n856), .Y(n469) );
NAND2X1 U421 ( .A(n443), .B(n442), .Y(n441) );
NOR2X1 U42200 ( .A(b_var[2]), .B(var_code[2]), .Y(n859) );
NOR2X1 U42201 ( .A(n281), .B(var_code[3]), .Y(n860) );
NOR2X1 U42202 ( .A(n859), .B(n859), .Y(n861) );
NOR2X1 U42203 ( .A(n860), .B(n860), .Y(n862) );
NAND2X1 U42204 ( .A(n861), .B(n862), .Y(n863) );
NAND2X1 U42205 ( .A(n863), .B(n863), .Y(n864) );
NAND2X1 U42206 ( .A(n864), .B(a_var[2]), .Y(n282) );
NAND2X1 U423 ( .A(b_var[2]), .B(b_var[2]), .Y(n281) );
NAND2X1 U42400 ( .A(n360), .B(cin), .Y(n865) );
NAND2X1 U42401 ( .A(n865), .B(n865), .Y(n866) );
NAND2X1 U42402 ( .A(n866), .B(n359), .Y(n867) );
NAND2X1 U42403 ( .A(n867), .B(n867), .Y(n868) );
NOR2X1 U42404 ( .A(n868), .B(n280), .Y(n443) );
NOR2X1 U42500 ( .A(b_var[0]), .B(n464), .Y(n869) );
NOR2X1 U42501 ( .A(n277), .B(n463), .Y(n870) );
NOR2X1 U42502 ( .A(n869), .B(n869), .Y(n871) );
NOR2X1 U42503 ( .A(n870), .B(n870), .Y(n872) );
NAND2X1 U42504 ( .A(n871), .B(n872), .Y(n873) );
NAND2X1 U42505 ( .A(n873), .B(n873), .Y(n874) );
NAND2X1 U42506 ( .A(n874), .B(a_var[0]), .Y(n275) );
NAND2X1 U426 ( .A(b_var[0]), .B(b_var[0]), .Y(n277) );
NOR2X1 U42700 ( .A(b_var[3]), .B(n464), .Y(n875) );
NOR2X1 U42701 ( .A(n272), .B(n463), .Y(n876) );
NOR2X1 U42702 ( .A(n875), .B(n875), .Y(n877) );
NOR2X1 U42703 ( .A(n876), .B(n876), .Y(n878) );
NAND2X1 U42704 ( .A(n877), .B(n878), .Y(n879) );
NAND2X1 U42705 ( .A(n879), .B(n879), .Y(n880) );
NAND2X1 U42706 ( .A(n880), .B(a_var[3]), .Y(n273) );
NAND2X1 U428 ( .A(b_var[3]), .B(b_var[3]), .Y(n272) );
NOR2X1 U42900 ( .A(b_var[4]), .B(n464), .Y(n881) );
NOR2X1 U42901 ( .A(n269), .B(n463), .Y(n882) );
NOR2X1 U42902 ( .A(n881), .B(n881), .Y(n883) );
NOR2X1 U42903 ( .A(n882), .B(n882), .Y(n884) );
NAND2X1 U42904 ( .A(n883), .B(n884), .Y(n885) );
NAND2X1 U42905 ( .A(n885), .B(n885), .Y(n886) );
NAND2X1 U42906 ( .A(n886), .B(a_var[4]), .Y(n270) );
NAND2X1 U430 ( .A(b_var[4]), .B(b_var[4]), .Y(n269) );
NAND2X1 U431 ( .A(a_var[5]), .B(a_var[5]), .Y(n265) );
NAND2X1 U432 ( .A(b_var[5]), .B(b_var[5]), .Y(n267) );
NAND2X1 U433 ( .A(a_var[6]), .B(a_var[6]), .Y(n262) );
NAND2X1 U434 ( .A(a_var[7]), .B(a_var[7]), .Y(n259) );
NAND2X1 U435 ( .A(b_var[7]), .B(b_var[7]), .Y(n286) );
NOR2X1 U43600 ( .A(b_var[8]), .B(n464), .Y(n887) );
NOR2X1 U43601 ( .A(n288), .B(n463), .Y(n888) );
NOR2X1 U43602 ( .A(n887), .B(n887), .Y(n889) );
NOR2X1 U43603 ( .A(n888), .B(n888), .Y(n890) );
NAND2X1 U43604 ( .A(n889), .B(n890), .Y(n891) );
NAND2X1 U43605 ( .A(n891), .B(n891), .Y(n892) );
NAND2X1 U43606 ( .A(n892), .B(a_var[8]), .Y(n256) );
NAND2X1 U437 ( .A(b_var[8]), .B(b_var[8]), .Y(n288) );
NOR2X1 U43800 ( .A(b_var[9]), .B(n464), .Y(n893) );
NOR2X1 U43801 ( .A(n253), .B(n463), .Y(n894) );
NOR2X1 U43802 ( .A(n893), .B(n893), .Y(n895) );
NOR2X1 U43803 ( .A(n894), .B(n894), .Y(n896) );
NAND2X1 U43804 ( .A(n895), .B(n896), .Y(n897) );
NAND2X1 U43805 ( .A(n897), .B(n897), .Y(n898) );
NAND2X1 U43806 ( .A(n898), .B(a_var[9]), .Y(n254) );
NAND2X1 U439 ( .A(b_var[9]), .B(b_var[9]), .Y(n253) );
NAND2X1 U440 ( .A(n300), .B(n300), .Y(n306) );
NAND2X1 U44100 ( .A(n303), .B(n303), .Y(n899) );
NAND2X1 U44101 ( .A(n493), .B(n493), .Y(n900) );
NAND2X1 U44102 ( .A(n899), .B(n900), .Y(n901) );
NOR2X1 U44103 ( .A(n902), .B(n302), .Y(n309) );
NAND2X1 U44104 ( .A(n901), .B(n901), .Y(n902) );
NAND2X1 U442 ( .A(n319), .B(n319), .Y(n322) );
NOR2X1 U44300 ( .A(b_var[14]), .B(n464), .Y(n903) );
NOR2X1 U44301 ( .A(n317), .B(n463), .Y(n904) );
NOR2X1 U44302 ( .A(n903), .B(n903), .Y(n905) );
NOR2X1 U44303 ( .A(n904), .B(n904), .Y(n906) );
NAND2X1 U44304 ( .A(n905), .B(n906), .Y(n907) );
NAND2X1 U44305 ( .A(n907), .B(n907), .Y(n908) );
NAND2X1 U44306 ( .A(n908), .B(a_var[14]), .Y(n313) );
NAND2X1 U444 ( .A(b_var[14]), .B(b_var[14]), .Y(n317) );
NOR2X1 U44500 ( .A(b_var[12]), .B(n464), .Y(n909) );
NOR2X1 U44501 ( .A(n304), .B(n463), .Y(n910) );
NOR2X1 U44502 ( .A(n909), .B(n909), .Y(n911) );
NOR2X1 U44503 ( .A(n910), .B(n910), .Y(n912) );
NAND2X1 U44504 ( .A(n911), .B(n912), .Y(n913) );
NAND2X1 U44505 ( .A(n913), .B(n913), .Y(n914) );
NAND2X1 U44506 ( .A(n914), .B(a_var[12]), .Y(n294) );
NAND2X1 U446 ( .A(b_var[12]), .B(b_var[12]), .Y(n304) );
NOR2X1 U44700 ( .A(b_var[13]), .B(n464), .Y(n915) );
NOR2X1 U44701 ( .A(n303), .B(n463), .Y(n916) );
NOR2X1 U44702 ( .A(n915), .B(n915), .Y(n917) );
NOR2X1 U44703 ( .A(n916), .B(n916), .Y(n918) );
NAND2X1 U44704 ( .A(n917), .B(n918), .Y(n919) );
NAND2X1 U44705 ( .A(n919), .B(n919), .Y(n920) );
NAND2X1 U44706 ( .A(n920), .B(a_var[13]), .Y(n298) );
NAND2X1 U448 ( .A(b_var[13]), .B(b_var[13]), .Y(n303) );
NOR2X1 U44900 ( .A(b_var[16]), .B(n464), .Y(n921) );
NOR2X1 U44901 ( .A(n331), .B(n463), .Y(n922) );
NOR2X1 U44902 ( .A(n921), .B(n921), .Y(n923) );
NOR2X1 U44903 ( .A(n922), .B(n922), .Y(n924) );
NAND2X1 U44904 ( .A(n923), .B(n924), .Y(n925) );
NAND2X1 U44905 ( .A(n925), .B(n925), .Y(n926) );
NAND2X1 U44906 ( .A(n926), .B(a_var[16]), .Y(n327) );
NAND2X1 U450 ( .A(b_var[16]), .B(b_var[16]), .Y(n331) );
NOR2X1 U45100 ( .A(b_var[17]), .B(n464), .Y(n927) );
NOR2X1 U45101 ( .A(n337), .B(n463), .Y(n928) );
NOR2X1 U45102 ( .A(n927), .B(n927), .Y(n929) );
NOR2X1 U45103 ( .A(n928), .B(n928), .Y(n930) );
NAND2X1 U45104 ( .A(n929), .B(n930), .Y(n931) );
NAND2X1 U45105 ( .A(n931), .B(n931), .Y(n932) );
NAND2X1 U45106 ( .A(n932), .B(a_var[17]), .Y(n329) );
NAND2X1 U452 ( .A(b_var[17]), .B(b_var[17]), .Y(n337) );
NAND2X1 U453 ( .A(anl), .B(b_var[18]), .Y(n355) );
NOR2X1 U45400 ( .A(b_var[18]), .B(var_code[2]), .Y(n933) );
NOR2X1 U45401 ( .A(n340), .B(var_code[3]), .Y(n934) );
NOR2X1 U45402 ( .A(n933), .B(n933), .Y(n935) );
NOR2X1 U45403 ( .A(n934), .B(n934), .Y(n936) );
NAND2X1 U45404 ( .A(n935), .B(n936), .Y(n937) );
NAND2X1 U45405 ( .A(n937), .B(n937), .Y(n938) );
NAND2X1 U45406 ( .A(n938), .B(a_var[18]), .Y(n341) );
NAND2X1 U455 ( .A(b_var[18]), .B(b_var[18]), .Y(n340) );
NAND2X1 U456 ( .A(a_var[19]), .B(a_var[19]), .Y(n346) );
NAND2X1 U457 ( .A(b_var[19]), .B(b_var[19]), .Y(n365) );
NAND2X1 U458 ( .A(a_var[20]), .B(a_var[20]), .Y(n362) );
NAND2X1 U459 ( .A(n399), .B(n399), .Y(n396) );
NAND2X1 U460 ( .A(n384), .B(n384), .Y(n379) );
NOR2X1 U46100 ( .A(b_var[22]), .B(var_code[2]), .Y(n939) );
NOR2X1 U46101 ( .A(n375), .B(var_code[3]), .Y(n940) );
NOR2X1 U46102 ( .A(n939), .B(n939), .Y(n941) );
NOR2X1 U46103 ( .A(n940), .B(n940), .Y(n942) );
NAND2X1 U46104 ( .A(n941), .B(n942), .Y(n943) );
NAND2X1 U46105 ( .A(n943), .B(n943), .Y(n944) );
NAND2X1 U46106 ( .A(n944), .B(a_var[22]), .Y(n376) );
NAND2X1 U462 ( .A(b_var[22]), .B(b_var[22]), .Y(n375) );
NAND2X1 U463 ( .A(a_var[21]), .B(a_var[21]), .Y(n370) );
NAND2X1 U464 ( .A(b_var[21]), .B(b_var[21]), .Y(n378) );
NAND2X1 U465 ( .A(a_var[23]), .B(a_var[23]), .Y(n386) );
NAND2X1 U466 ( .A(b_var[23]), .B(b_var[23]), .Y(n393) );
NOR2X1 U46700 ( .A(b_var[24]), .B(n464), .Y(n945) );
NOR2X1 U46701 ( .A(n390), .B(n463), .Y(n946) );
NOR2X1 U46702 ( .A(n945), .B(n945), .Y(n947) );
NOR2X1 U46703 ( .A(n946), .B(n946), .Y(n948) );
NAND2X1 U46704 ( .A(n947), .B(n948), .Y(n949) );
NAND2X1 U46705 ( .A(n949), .B(n949), .Y(n950) );
NAND2X1 U46706 ( .A(n950), .B(a_var[24]), .Y(n391) );
NAND2X1 U468 ( .A(b_var[24]), .B(b_var[24]), .Y(n390) );
NOR2X1 U46900 ( .A(b_var[25]), .B(n464), .Y(n951) );
NOR2X1 U46901 ( .A(n411), .B(n463), .Y(n952) );
NOR2X1 U46902 ( .A(n951), .B(n951), .Y(n953) );
NOR2X1 U46903 ( .A(n952), .B(n952), .Y(n954) );
NAND2X1 U46904 ( .A(n953), .B(n954), .Y(n955) );
NAND2X1 U46905 ( .A(n955), .B(n955), .Y(n956) );
NAND2X1 U46906 ( .A(n956), .B(a_var[25]), .Y(n401) );
NAND2X1 U470 ( .A(b_var[25]), .B(b_var[25]), .Y(n411) );
NAND2X1 U471 ( .A(a_var[27]), .B(a_var[27]), .Y(n419) );
NAND2X1 U472 ( .A(b_var[27]), .B(b_var[27]), .Y(n427) );
NOR2X1 U47300 ( .A(b_var[28]), .B(n464), .Y(n957) );
NOR2X1 U47301 ( .A(n433), .B(n463), .Y(n958) );
NOR2X1 U47302 ( .A(n957), .B(n957), .Y(n959) );
NOR2X1 U47303 ( .A(n958), .B(n958), .Y(n960) );
NAND2X1 U47304 ( .A(n959), .B(n960), .Y(n961) );
NAND2X1 U47305 ( .A(n961), .B(n961), .Y(n962) );
NAND2X1 U47306 ( .A(n962), .B(a_var[28]), .Y(n425) );
NAND2X1 U474 ( .A(b_var[28]), .B(b_var[28]), .Y(n433) );
NAND2X1 U475 ( .A(anl), .B(b_var[29]), .Y(n454) );
NOR2X1 U47600 ( .A(b_var[29]), .B(var_code[2]), .Y(n963) );
NOR2X1 U47601 ( .A(n436), .B(var_code[3]), .Y(n964) );
NOR2X1 U47602 ( .A(n963), .B(n963), .Y(n965) );
NOR2X1 U47603 ( .A(n964), .B(n964), .Y(n966) );
NAND2X1 U47604 ( .A(n965), .B(n966), .Y(n967) );
NAND2X1 U47605 ( .A(n967), .B(n967), .Y(n968) );
NAND2X1 U47606 ( .A(n968), .B(a_var[29]), .Y(n437) );
NAND2X1 U477 ( .A(b_var[29]), .B(b_var[29]), .Y(n436) );
NAND2X1 U478 ( .A(a_var[30]), .B(a_var[30]), .Y(n445) );
NAND2X1 U479 ( .A(b_var[6]), .B(b_var[6]), .Y(n285) );
NAND2X1 U480 ( .A(b_var[20]), .B(b_var[20]), .Y(n373) );
NAND2X1 U481 ( .A(b_var[30]), .B(b_var[30]), .Y(n459) );
NOR2X1 U48200 ( .A(b_var[9]), .B(n462), .Y(n969) );
NOR2X1 U48201 ( .A(n253), .B(n461), .Y(n970) );
NOR2X1 U48202 ( .A(n969), .B(n969), .Y(n971) );
NOR2X1 U48203 ( .A(n970), .B(n970), .Y(n972) );
NAND2X1 U48204 ( .A(n971), .B(n972), .Y(n255) );
NOR2X1 U48300 ( .A(b_var[6]), .B(n462), .Y(n973) );
NOR2X1 U48301 ( .A(n285), .B(n461), .Y(n974) );
NOR2X1 U48302 ( .A(n973), .B(n973), .Y(n975) );
NOR2X1 U48303 ( .A(n974), .B(n974), .Y(n976) );
NAND2X1 U48304 ( .A(n975), .B(n976), .Y(n263) );
NOR2X1 U48400 ( .A(b_var[6]), .B(n464), .Y(n977) );
NOR2X1 U48401 ( .A(n285), .B(n463), .Y(n978) );
NOR2X1 U48402 ( .A(n977), .B(n977), .Y(n979) );
NOR2X1 U48403 ( .A(n978), .B(n978), .Y(n980) );
NAND2X1 U48404 ( .A(n979), .B(n980), .Y(n261) );
NOR2X1 U48500 ( .A(b_var[5]), .B(var_code[0]), .Y(n981) );
NOR2X1 U48501 ( .A(n267), .B(var_code[1]), .Y(n982) );
NOR2X1 U48502 ( .A(n981), .B(n981), .Y(n983) );
NOR2X1 U48503 ( .A(n982), .B(n982), .Y(n984) );
NAND2X1 U48504 ( .A(n983), .B(n984), .Y(n266) );
NOR2X1 U48600 ( .A(b_var[5]), .B(var_code[2]), .Y(n985) );
NOR2X1 U48601 ( .A(n267), .B(var_code[3]), .Y(n986) );
NOR2X1 U48602 ( .A(n985), .B(n985), .Y(n987) );
NOR2X1 U48603 ( .A(n986), .B(n986), .Y(n988) );
NAND2X1 U48604 ( .A(n987), .B(n988), .Y(n264) );
NOR2X1 U487 ( .A(n493), .B(n267), .Y(n268) );
NOR2X1 U48800 ( .A(n284), .B(n477), .Y(n989) );
NOR2X1 U48801 ( .A(n989), .B(n989), .Y(n990) );
NOR2X1 U48802 ( .A(n990), .B(n268), .Y(n474) );
NOR2X1 U48900 ( .A(b_var[4]), .B(n462), .Y(n991) );
NOR2X1 U48901 ( .A(n269), .B(n461), .Y(n992) );
NOR2X1 U48902 ( .A(n991), .B(n991), .Y(n993) );
NOR2X1 U48903 ( .A(n992), .B(n992), .Y(n994) );
NAND2X1 U48904 ( .A(n993), .B(n994), .Y(n271) );
NOR2X1 U49000 ( .A(b_var[3]), .B(n462), .Y(n995) );
NOR2X1 U49001 ( .A(n272), .B(n461), .Y(n996) );
NOR2X1 U49002 ( .A(n995), .B(n995), .Y(n997) );
NOR2X1 U49003 ( .A(n996), .B(n996), .Y(n998) );
NAND2X1 U49004 ( .A(n997), .B(n998), .Y(n274) );
NOR2X1 U49100 ( .A(b_var[0]), .B(n462), .Y(n999) );
NOR2X1 U49101 ( .A(n277), .B(n461), .Y(n1000) );
NOR2X1 U49102 ( .A(n999), .B(n999), .Y(n1001) );
NOR2X1 U49103 ( .A(n1000), .B(n1000), .Y(n1002) );
NAND2X1 U49104 ( .A(n1001), .B(n1002), .Y(n276) );
NOR2X1 U49200 ( .A(b_var[1]), .B(n360), .Y(n1003) );
NOR2X1 U49201 ( .A(n1003), .B(n1003), .Y(n1004) );
NAND2X1 U49202 ( .A(n1004), .B(n278), .Y(n279) );
NOR2X1 U493 ( .A(n493), .B(n279), .Y(n280) );
NOR2X1 U49400 ( .A(b_var[2]), .B(var_code[0]), .Y(n1005) );
NOR2X1 U49401 ( .A(n281), .B(var_code[1]), .Y(n1006) );
NOR2X1 U49402 ( .A(n1005), .B(n1005), .Y(n1007) );
NOR2X1 U49403 ( .A(n1006), .B(n1006), .Y(n1008) );
NAND2X1 U49404 ( .A(n1007), .B(n1008), .Y(n283) );
NOR2X1 U495 ( .A(n469), .B(n468), .Y(n467) );
NOR2X1 U496 ( .A(n472), .B(n471), .Y(n470) );
NOR2X1 U497 ( .A(n474), .B(n475), .Y(n484) );
NAND2X1 U49800 ( .A(b_var[5]), .B(anl), .Y(n1009) );
NAND2X1 U49801 ( .A(n1009), .B(n1009), .Y(n1010) );
NAND2X1 U49802 ( .A(n1010), .B(n473), .Y(n481) );
NOR2X1 U49900 ( .A(n288), .B(n493), .Y(n1011) );
NOR2X1 U49901 ( .A(n1011), .B(n1011), .Y(n1012) );
NAND2X1 U49902 ( .A(n1012), .B(n486), .Y(n289) );
NOR2X1 U50000 ( .A(n486), .B(cout7), .Y(n1013) );
NOR2X1 U50001 ( .A(n1013), .B(n1013), .Y(n1014) );
NAND2X1 U50002 ( .A(n1014), .B(n289), .Y(n489) );
NOR2X1 U501 ( .A(n489), .B(n488), .Y(n487) );
NOR2X1 U50200 ( .A(n296), .B(n293), .Y(n1015) );
NOR2X1 U50201 ( .A(n1015), .B(n1015), .Y(n1016) );
NAND2X1 U50202 ( .A(n1016), .B(n297), .Y(result[11]) );
NAND2X1 U50300 ( .A(b_var[12]), .B(anl), .Y(n1017) );
NAND2X1 U50301 ( .A(n1017), .B(n1017), .Y(n1018) );
NAND2X1 U50302 ( .A(n1018), .B(n300), .Y(n311) );
NOR2X1 U50400 ( .A(n300), .B(n307), .Y(n1019) );
NOR2X1 U50401 ( .A(n1019), .B(n1019), .Y(n1020) );
NAND2X1 U50402 ( .A(n1020), .B(n311), .Y(n301) );
NAND2X1 U50500 ( .A(n301), .B(n302), .Y(n1021) );
NAND2X1 U50501 ( .A(n1021), .B(n1021), .Y(n1025) );
NAND2X1 U50502 ( .A(n301), .B(n301), .Y(n1022) );
NAND2X1 U50503 ( .A(n1022), .B(n312), .Y(n1023) );
NAND2X1 U50504 ( .A(n1023), .B(n1023), .Y(n1024) );
NOR2X1 U50505 ( .A(n1024), .B(n1025), .Y(result[13]) );
NOR2X1 U506 ( .A(n493), .B(n304), .Y(n305) );
NOR2X1 U50700 ( .A(n306), .B(n305), .Y(n1026) );
NOR2X1 U50701 ( .A(n1026), .B(n1026), .Y(n1027) );
NOR2X1 U50702 ( .A(n1027), .B(n312), .Y(n308) );
NAND2X1 U50800 ( .A(n312), .B(anl), .Y(n1028) );
NAND2X1 U50801 ( .A(n1028), .B(n1028), .Y(n1029) );
NAND2X1 U50802 ( .A(n1029), .B(b_var[13]), .Y(n310) );
NOR2X1 U50900 ( .A(n312), .B(n311), .Y(n1030) );
NOR2X1 U50901 ( .A(n1030), .B(n1030), .Y(n1031) );
NAND2X1 U50902 ( .A(n1031), .B(n310), .Y(n320) );
NOR2X1 U510 ( .A(n321), .B(n320), .Y(n316) );
NOR2X1 U51100 ( .A(n316), .B(n322), .Y(n1032) );
NOR2X1 U51101 ( .A(n1032), .B(n1032), .Y(n1033) );
NAND2X1 U51102 ( .A(n1033), .B(n315), .Y(result[14]) );
NOR2X1 U51200 ( .A(n493), .B(n317), .Y(n1034) );
NOR2X1 U51201 ( .A(n1034), .B(n1034), .Y(n1035) );
NAND2X1 U51202 ( .A(n1035), .B(n319), .Y(n318) );
NOR2X1 U513 ( .A(n326), .B(n323), .Y(n335) );
NAND2X1 U51400 ( .A(n326), .B(b_var[15]), .Y(n1036) );
NAND2X1 U51401 ( .A(n1036), .B(n1036), .Y(n1037) );
NAND2X1 U51402 ( .A(n1037), .B(anl), .Y(n324) );
NOR2X1 U51500 ( .A(b_var[16]), .B(n462), .Y(n1038) );
NOR2X1 U51501 ( .A(n331), .B(n461), .Y(n1039) );
NOR2X1 U51502 ( .A(n1038), .B(n1038), .Y(n1040) );
NOR2X1 U51503 ( .A(n1039), .B(n1039), .Y(n1041) );
NAND2X1 U51504 ( .A(n1040), .B(n1041), .Y(n328) );
NOR2X1 U51600 ( .A(b_var[17]), .B(n462), .Y(n1042) );
NOR2X1 U51601 ( .A(n337), .B(n461), .Y(n1043) );
NOR2X1 U51602 ( .A(n1042), .B(n1042), .Y(n1044) );
NOR2X1 U51603 ( .A(n1043), .B(n1043), .Y(n1045) );
NAND2X1 U51604 ( .A(n1044), .B(n1045), .Y(n330) );
NOR2X1 U51700 ( .A(n331), .B(n493), .Y(n1046) );
NOR2X1 U51701 ( .A(n1046), .B(n1046), .Y(n1047) );
NAND2X1 U51702 ( .A(n1047), .B(n333), .Y(n334) );
NOR2X1 U51800 ( .A(n333), .B(n332), .Y(n1048) );
NOR2X1 U51801 ( .A(n1048), .B(n1048), .Y(n1049) );
NAND2X1 U51802 ( .A(n1049), .B(n334), .Y(n349) );
NAND2X1 U51900 ( .A(n336), .B(n349), .Y(n1050) );
NAND2X1 U51901 ( .A(n1050), .B(n1050), .Y(n1051) );
NAND2X1 U51902 ( .A(n1051), .B(n350), .Y(n339) );
NOR2X1 U52000 ( .A(n337), .B(n493), .Y(n1052) );
NOR2X1 U52001 ( .A(n1052), .B(n1052), .Y(n1053) );
NAND2X1 U52002 ( .A(n1053), .B(n351), .Y(n338) );
NOR2X1 U52100 ( .A(b_var[18]), .B(var_code[0]), .Y(n1054) );
NOR2X1 U52101 ( .A(n340), .B(var_code[1]), .Y(n1055) );
NOR2X1 U52102 ( .A(n1054), .B(n1054), .Y(n1056) );
NOR2X1 U52103 ( .A(n1055), .B(n1055), .Y(n1057) );
NAND2X1 U52104 ( .A(n1056), .B(n1057), .Y(n342) );
NOR2X1 U52200 ( .A(b_var[19]), .B(var_code[0]), .Y(n1058) );
NOR2X1 U52201 ( .A(n365), .B(var_code[1]), .Y(n1059) );
NOR2X1 U52202 ( .A(n1058), .B(n1058), .Y(n1060) );
NOR2X1 U52203 ( .A(n1059), .B(n1059), .Y(n1061) );
NAND2X1 U52204 ( .A(n1060), .B(n1061), .Y(n347) );
NOR2X1 U52300 ( .A(b_var[19]), .B(var_code[2]), .Y(n1062) );
NOR2X1 U52301 ( .A(n365), .B(var_code[3]), .Y(n1063) );
NOR2X1 U52302 ( .A(n1062), .B(n1062), .Y(n1064) );
NOR2X1 U52303 ( .A(n1063), .B(n1063), .Y(n1065) );
NAND2X1 U52304 ( .A(n1064), .B(n1065), .Y(n345) );
NAND2X1 U52400 ( .A(n351), .B(anl), .Y(n1066) );
NAND2X1 U52401 ( .A(n1066), .B(n1066), .Y(n1067) );
NAND2X1 U52402 ( .A(n1067), .B(b_var[17]), .Y(n348) );
NOR2X1 U52500 ( .A(n351), .B(n349), .Y(n1068) );
NOR2X1 U52501 ( .A(n1068), .B(n1068), .Y(n1069) );
NAND2X1 U52502 ( .A(n1069), .B(n348), .Y(n353) );
NOR2X1 U526 ( .A(n351), .B(n350), .Y(n352) );
NOR2X1 U52700 ( .A(n353), .B(n352), .Y(n1070) );
NOR2X1 U52701 ( .A(n1070), .B(n1070), .Y(n1071) );
NAND2X1 U52702 ( .A(n1071), .B(n356), .Y(n354) );
NOR2X1 U52800 ( .A(n356), .B(n355), .Y(n1072) );
NOR2X1 U52801 ( .A(n1072), .B(n1072), .Y(n1073) );
NAND2X1 U52802 ( .A(n1073), .B(n354), .Y(n357) );
NOR2X1 U52900 ( .A(n366), .B(n357), .Y(n1074) );
NOR2X1 U52901 ( .A(n1074), .B(n1074), .Y(n1075) );
NAND2X1 U52902 ( .A(n1075), .B(n364), .Y(n358) );
NOR2X1 U53000 ( .A(b_var[20]), .B(var_code[0]), .Y(n1076) );
NOR2X1 U53001 ( .A(n373), .B(var_code[1]), .Y(n1077) );
NOR2X1 U53002 ( .A(n1076), .B(n1076), .Y(n1078) );
NOR2X1 U53003 ( .A(n1077), .B(n1077), .Y(n1079) );
NAND2X1 U53004 ( .A(n1078), .B(n1079), .Y(n363) );
NOR2X1 U53100 ( .A(b_var[20]), .B(var_code[2]), .Y(n1080) );
NOR2X1 U53101 ( .A(n373), .B(var_code[3]), .Y(n1081) );
NOR2X1 U53102 ( .A(n1080), .B(n1080), .Y(n1082) );
NOR2X1 U53103 ( .A(n1081), .B(n1081), .Y(n1083) );
NAND2X1 U53104 ( .A(n1082), .B(n1083), .Y(n361) );
NOR2X1 U53200 ( .A(n374), .B(n367), .Y(n1084) );
NOR2X1 U53201 ( .A(n1084), .B(n1084), .Y(n1085) );
NAND2X1 U53202 ( .A(n1085), .B(n372), .Y(n368) );
NOR2X1 U53300 ( .A(b_var[21]), .B(var_code[0]), .Y(n1086) );
NOR2X1 U53301 ( .A(n378), .B(var_code[1]), .Y(n1087) );
NOR2X1 U53302 ( .A(n1086), .B(n1086), .Y(n1088) );
NOR2X1 U53303 ( .A(n1087), .B(n1087), .Y(n1089) );
NAND2X1 U53304 ( .A(n1088), .B(n1089), .Y(n371) );
NOR2X1 U53400 ( .A(b_var[21]), .B(var_code[2]), .Y(n1090) );
NOR2X1 U53401 ( .A(n378), .B(var_code[3]), .Y(n1091) );
NOR2X1 U53402 ( .A(n1090), .B(n1090), .Y(n1092) );
NOR2X1 U53403 ( .A(n1091), .B(n1091), .Y(n1093) );
NAND2X1 U53404 ( .A(n1092), .B(n1093), .Y(n369) );
NOR2X1 U53500 ( .A(n384), .B(n400), .Y(n1094) );
NOR2X1 U53501 ( .A(n379), .B(n409), .Y(n1095) );
NOR2X1 U53502 ( .A(n1094), .B(n1094), .Y(n1096) );
NOR2X1 U53503 ( .A(n1095), .B(n1095), .Y(n1097) );
NAND2X1 U53504 ( .A(n1096), .B(n1097), .Y(result[21]) );
NAND2X1 U53600 ( .A(n380), .B(n383), .Y(n1098) );
NAND2X1 U53601 ( .A(n1098), .B(n1098), .Y(n1102) );
NAND2X1 U53602 ( .A(n380), .B(n380), .Y(n1099) );
NAND2X1 U53603 ( .A(n1099), .B(n382), .Y(n1100) );
NAND2X1 U53604 ( .A(n1100), .B(n1100), .Y(n1101) );
NOR2X1 U53605 ( .A(n1101), .B(n1102), .Y(result[22]) );
NAND2X1 U53700 ( .A(anl), .B(b_var[22]), .Y(n1103) );
NAND2X1 U53701 ( .A(n1103), .B(n1103), .Y(n1104) );
NAND2X1 U53702 ( .A(n1104), .B(n383), .Y(n395) );
NOR2X1 U53800 ( .A(n384), .B(n394), .Y(n1105) );
NOR2X1 U53801 ( .A(n1105), .B(n1105), .Y(n1106) );
NAND2X1 U53802 ( .A(n1106), .B(n395), .Y(n398) );
NOR2X1 U53900 ( .A(b_var[23]), .B(n462), .Y(n1107) );
NOR2X1 U53901 ( .A(n393), .B(n461), .Y(n1108) );
NOR2X1 U53902 ( .A(n1107), .B(n1107), .Y(n1109) );
NOR2X1 U53903 ( .A(n1108), .B(n1108), .Y(n1110) );
NAND2X1 U53904 ( .A(n1109), .B(n1110), .Y(n387) );
NOR2X1 U54000 ( .A(b_var[23]), .B(n464), .Y(n1111) );
NOR2X1 U54001 ( .A(n393), .B(n463), .Y(n1112) );
NOR2X1 U54002 ( .A(n1111), .B(n1111), .Y(n1113) );
NOR2X1 U54003 ( .A(n1112), .B(n1112), .Y(n1114) );
NAND2X1 U54004 ( .A(n1113), .B(n1114), .Y(n385) );
NOR2X1 U54100 ( .A(n493), .B(n393), .Y(n1115) );
NOR2X1 U54101 ( .A(n1115), .B(n1115), .Y(n1116) );
NAND2X1 U54102 ( .A(n1116), .B(n399), .Y(n397) );
NOR2X1 U54200 ( .A(n399), .B(n398), .Y(n1117) );
NOR2X1 U54201 ( .A(n1117), .B(n1117), .Y(n1118) );
NAND2X1 U54202 ( .A(n1118), .B(n397), .Y(n405) );
NAND2X1 U54300 ( .A(n406), .B(b_var[24]), .Y(n1119) );
NAND2X1 U54301 ( .A(n1119), .B(n1119), .Y(n1120) );
NAND2X1 U54302 ( .A(n1120), .B(anl), .Y(n404) );
NOR2X1 U54400 ( .A(n406), .B(n403), .Y(n1121) );
NOR2X1 U54401 ( .A(n1121), .B(n1121), .Y(n1122) );
NAND2X1 U54402 ( .A(n1122), .B(n404), .Y(n410) );
NOR2X1 U54500 ( .A(n406), .B(n405), .Y(n1123) );
NOR2X1 U54501 ( .A(n1123), .B(n1123), .Y(n1124) );
NAND2X1 U54502 ( .A(n1124), .B(n404), .Y(n413) );
NAND2X1 U54600 ( .A(n407), .B(n414), .Y(n1125) );
NAND2X1 U54601 ( .A(n1125), .B(n1125), .Y(n1129) );
NAND2X1 U54602 ( .A(n407), .B(n407), .Y(n1126) );
NAND2X1 U54603 ( .A(n1126), .B(n408), .Y(n1127) );
NAND2X1 U54604 ( .A(n1127), .B(n1127), .Y(n1128) );
NOR2X1 U54605 ( .A(n1128), .B(n1129), .Y(result[25]) );
NOR2X1 U54700 ( .A(n493), .B(n411), .Y(n1130) );
NOR2X1 U54701 ( .A(n1130), .B(n1130), .Y(n1131) );
NAND2X1 U54702 ( .A(n1131), .B(n414), .Y(n412) );
NOR2X1 U54800 ( .A(n414), .B(n413), .Y(n1132) );
NOR2X1 U54801 ( .A(n1132), .B(n1132), .Y(n1133) );
NAND2X1 U54802 ( .A(n1133), .B(n412), .Y(n422) );
NOR2X1 U54900 ( .A(n416), .B(n423), .Y(n1134) );
NOR2X1 U54901 ( .A(n1134), .B(n1134), .Y(n1135) );
NAND2X1 U54902 ( .A(n1135), .B(n415), .Y(result[26]) );
NOR2X1 U550 ( .A(n423), .B(n417), .Y(n431) );
NOR2X1 U55100 ( .A(b_var[27]), .B(n462), .Y(n1136) );
NOR2X1 U55101 ( .A(n427), .B(n461), .Y(n1137) );
NOR2X1 U55102 ( .A(n1136), .B(n1136), .Y(n1138) );
NOR2X1 U55103 ( .A(n1137), .B(n1137), .Y(n1139) );
NAND2X1 U55104 ( .A(n1138), .B(n1139), .Y(n420) );
NOR2X1 U55200 ( .A(b_var[27]), .B(n464), .Y(n1140) );
NOR2X1 U55201 ( .A(n427), .B(n463), .Y(n1141) );
NOR2X1 U55202 ( .A(n1140), .B(n1140), .Y(n1142) );
NOR2X1 U55203 ( .A(n1141), .B(n1141), .Y(n1143) );
NAND2X1 U55204 ( .A(n1142), .B(n1143), .Y(n418) );
NAND2X1 U55300 ( .A(n423), .B(b_var[26]), .Y(n1144) );
NAND2X1 U55301 ( .A(n1144), .B(n1144), .Y(n1145) );
NAND2X1 U55302 ( .A(n1145), .B(anl), .Y(n421) );
NOR2X1 U55400 ( .A(n431), .B(n428), .Y(n1146) );
NOR2X1 U55401 ( .A(n1146), .B(n1146), .Y(n1147) );
NAND2X1 U55402 ( .A(n1147), .B(n429), .Y(n424) );
NOR2X1 U55500 ( .A(b_var[28]), .B(n462), .Y(n1148) );
NOR2X1 U55501 ( .A(n433), .B(n461), .Y(n1149) );
NOR2X1 U55502 ( .A(n1148), .B(n1148), .Y(n1150) );
NOR2X1 U55503 ( .A(n1149), .B(n1149), .Y(n1151) );
NAND2X1 U55504 ( .A(n1150), .B(n1151), .Y(n426) );
NOR2X1 U55600 ( .A(n493), .B(n427), .Y(n1152) );
NOR2X1 U55601 ( .A(n1152), .B(n1152), .Y(n1153) );
NAND2X1 U55602 ( .A(n1153), .B(n429), .Y(n430) );
NOR2X1 U55700 ( .A(n429), .B(n428), .Y(n1154) );
NOR2X1 U55701 ( .A(n1154), .B(n1154), .Y(n1155) );
NAND2X1 U55702 ( .A(n1155), .B(n430), .Y(n448) );
NAND2X1 U55800 ( .A(n432), .B(n448), .Y(n1156) );
NAND2X1 U55801 ( .A(n1156), .B(n1156), .Y(n1157) );
NAND2X1 U55802 ( .A(n1157), .B(n449), .Y(n435) );
NOR2X1 U55900 ( .A(n433), .B(n493), .Y(n1158) );
NOR2X1 U55901 ( .A(n1158), .B(n1158), .Y(n1159) );
NAND2X1 U55902 ( .A(n1159), .B(n450), .Y(n434) );
NOR2X1 U56000 ( .A(b_var[29]), .B(var_code[0]), .Y(n1160) );
NOR2X1 U56001 ( .A(n436), .B(var_code[1]), .Y(n1161) );
NOR2X1 U56002 ( .A(n1160), .B(n1160), .Y(n1162) );
NOR2X1 U56003 ( .A(n1161), .B(n1161), .Y(n1163) );
NAND2X1 U56004 ( .A(n1162), .B(n1163), .Y(n438) );
NOR2X1 U56100 ( .A(b_var[30]), .B(var_code[0]), .Y(n1164) );
NOR2X1 U56101 ( .A(n459), .B(var_code[1]), .Y(n1165) );
NOR2X1 U56102 ( .A(n1164), .B(n1164), .Y(n1166) );
NOR2X1 U56103 ( .A(n1165), .B(n1165), .Y(n1167) );
NAND2X1 U56104 ( .A(n1166), .B(n1167), .Y(n446) );
NOR2X1 U56200 ( .A(b_var[30]), .B(var_code[2]), .Y(n1168) );
NOR2X1 U56201 ( .A(n459), .B(var_code[3]), .Y(n1169) );
NOR2X1 U56202 ( .A(n1168), .B(n1168), .Y(n1170) );
NOR2X1 U56203 ( .A(n1169), .B(n1169), .Y(n1171) );
NAND2X1 U56204 ( .A(n1170), .B(n1171), .Y(n444) );
NAND2X1 U56300 ( .A(n450), .B(anl), .Y(n1172) );
NAND2X1 U56301 ( .A(n1172), .B(n1172), .Y(n1173) );
NAND2X1 U56302 ( .A(n1173), .B(b_var[28]), .Y(n447) );
NOR2X1 U56400 ( .A(n450), .B(n448), .Y(n1174) );
NOR2X1 U56401 ( .A(n1174), .B(n1174), .Y(n1175) );
NAND2X1 U56402 ( .A(n1175), .B(n447), .Y(n452) );
NOR2X1 U565 ( .A(n450), .B(n449), .Y(n451) );
NOR2X1 U56600 ( .A(n452), .B(n451), .Y(n1176) );
NOR2X1 U56601 ( .A(n1176), .B(n1176), .Y(n1177) );
NAND2X1 U56602 ( .A(n1177), .B(n455), .Y(n453) );
NOR2X1 U56700 ( .A(n460), .B(n456), .Y(n1178) );
NOR2X1 U56701 ( .A(n1178), .B(n1178), .Y(n1179) );
NAND2X1 U56702 ( .A(n1179), .B(n458), .Y(n457) );
NOR2X1 U56800 ( .A(b_var[31]), .B(n462), .Y(n1180) );
NOR2X1 U56801 ( .A(n492), .B(n461), .Y(n1181) );
NOR2X1 U56802 ( .A(n1180), .B(n1180), .Y(n1182) );
NOR2X1 U56803 ( .A(n1181), .B(n1181), .Y(n1183) );
NAND2X1 U56804 ( .A(n1182), .B(n1183), .Y(n466) );
NAND2X1 U56900 ( .A(n494), .B(cout30), .Y(n1184) );
NAND2X1 U56901 ( .A(n1184), .B(n1184), .Y(n1188) );
NAND2X1 U56902 ( .A(n494), .B(n494), .Y(n1185) );
NAND2X1 U56903 ( .A(n1185), .B(n491), .Y(n1186) );
NAND2X1 U56904 ( .A(n1186), .B(n1186), .Y(n1187) );
NOR2X1 U56905 ( .A(n1187), .B(n1188), .Y(result[31]) );
NOR2X1 U57000 ( .A(n477), .B(n475), .Y(n1189) );
NOR2X1 U57001 ( .A(n473), .B(n476), .Y(n1190) );
NOR2X1 U57002 ( .A(n1189), .B(n1189), .Y(n1191) );
NOR2X1 U57003 ( .A(n1190), .B(n1190), .Y(n1192) );
NAND2X1 U57004 ( .A(n1191), .B(n1192), .Y(result[5]) );
endmodule